module sink2 (clk, reset, req, ack, data);

	parameter id = 0;

	input clk, reset, req;

	input [`SIZE-1:0] data;

	output reg ack;

	reg req_old;

	always @(posedge clk or posedge reset) begin

		if (reset) begin

			req_old <= 0;

			ack <= 0;

		end else begin

			req_old <= req;

			if (req ^ req_old) begin

				$display("[%g] sink %g: received %g", $time, id, data);

				ack <= ~ack;

			end

		end
	end

endmodule
